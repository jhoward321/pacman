module maze (input [5:0] x_tile, y_tile, output up, down, left, right);
//takes in current sprite x and y tiles, outputs which directions sprite can move next

//need to convert 639x479 to 28x36 tiles

//how do I set each block to traversable or not? might be easier in c

